----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:00:17 03/04/2015 
-- Design Name: 
-- Module Name:    INST_MEM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity INST_MEM is
PORT( INST_ADDR: in STD_LOGIC;
		INST_IN: in STD_LOGIC_VECTOR (15 downto 0);
		INST_OUT: out STD_LOGIC_VECTOR (15 downto 0));
		
end INST_MEM;

architecture Behavioral of INST_MEM is

begin


end Behavioral;

